-- arm_one_nios.vhd

-- Generated using ACDS version 17.0 595

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity arm_one_nios_main is
	port (
	
		----------FPGA connections-------------
		CLOCK_50						: in std_logic;
		
		LEDR							: out std_logic_vector(9 downto 0);
		
		SDRAM_ADDR					: out std_logic_vector(10 downto 0);
		SDRAM_BA						: out std_logic_vector(1 downto 0);
		SDRAM_CAS_N					: out std_logic;
		SDRAM_CKE					: out std_logic;
		SDRAM_CS_N					: out std_logic;
		SDRAM_DQ						: inout std_logic_vector(15 downto 0);
		SDRAM_DQM					: out std_logic_vector(1 downto 0);
		SDRAM_RAS_N					: out std_logic;
		SDRAM_WE_N					: out std_logic;
		
		----------HPS connections--------------
		HPS_CONV_USB				: inout std_logic;
		
		HPS_DDR3_ADDR				: out std_logic_vector(14 downto 0);
		HPS_DDR3_BA					: out std_logic_vector(2 downto 0);
		HPS_DDR3_CAS_N				: out std_logic;
		HPS_DDR3_CKE				: out std_logic;
		HPS_DDR3_CK_N				: out std_logic;
		HPS_DDR3_CK_P				: out std_logic;
		HPS_DDR3_CS_N				: out std_logic;
		HPS_DDR3_DM					: out std_logic_vector(3 downto 0);
		HPS_DDR3_DQ					: inout std_logic_vector(31 downto 0);
		HPS_DDR3_DQS_N				: inout std_logic_vector(3 downto 0);
		HPS_DDR3_DQS_P				: inout std_logic_vector(3 downto 0);
		HPS_DDR3_ODT				: out std_logic;
		HPS_DDR3_RAS_N				: out std_logic;
		HPS_DDR3_RESET_N			: out std_logic;
		HPS_DDR3_RZQ				: in std_logic;
		HPS_DDR3_WE_N				: out std_logic;
		
		HPS_ENET_TX_CLK			: out std_logic;
		HPS_ENET_TX_EN				: out std_logic;
		HPS_ENET_TX_DATA			: out std_logic_vector(3 downto 0);
		HPS_ENET_RX_CLK			: in std_logic;
		HPS_ENET_RX_DV				: in std_logic;
		HPS_ENET_RX_DATA			: in std_logic_vector(3 downto 0);
		HPS_ENET_MDIO				: inout std_logic;
		HPS_ENET_MDC				: out std_logic;
		HPS_ENET_INT_N				: inout std_logic;

		HPS_KEY						: inout std_logic;
		
		HPS_SD_CLK					: out std_logic;
		HPS_SD_CMD					: inout std_logic;
		HPS_SD_DATA					: inout std_logic_vector(3 downto 0);
		
		HPS_UART_RX					: in std_logic;
		HPS_UART_TX					: out std_logic;
		
		HPS_USB_CLKOUT				: in std_logic;
		HPS_USB_DATA				: inout std_logic_vector(7 downto 0);
		HPS_USB_DIR					: in std_logic;
		HPS_USB_NXT					: in std_logic;
		HPS_USB_STP					: out std_logic
	);
end arm_one_nios_main;

architecture main of arm_one_nios_main is
	component arm_one_nios is
		port (
			clk_clk										: in std_logic;
			reset_reset_n								: in std_logic;
			
			hps_0_h2f_reset_reset_n					: out std_logic;
			
			hps_io_hps_io_emac1_inst_TX_CLK		: out std_logic;
			hps_io_hps_io_emac1_inst_TX_CTL		: out std_logic;
			hps_io_hps_io_emac1_inst_TXD0			: out std_logic;
			hps_io_hps_io_emac1_inst_TXD1			: out std_logic;
			hps_io_hps_io_emac1_inst_TXD2			: out std_logic;
			hps_io_hps_io_emac1_inst_TXD3			: out std_logic;
			hps_io_hps_io_emac1_inst_RX_CLK		: in std_logic;
			hps_io_hps_io_emac1_inst_RX_CTL		: in std_logic;
			hps_io_hps_io_emac1_inst_RXD0			: in std_logic;
			hps_io_hps_io_emac1_inst_RXD1			: in std_logic;
			hps_io_hps_io_emac1_inst_RXD2			: in std_logic;
			hps_io_hps_io_emac1_inst_RXD3			: in std_logic;
			hps_io_hps_io_emac1_inst_MDIO			: inout std_logic;
			hps_io_hps_io_emac1_inst_MDC			: out std_logic;
			
			hps_io_hps_io_sdio_inst_CLK			: out std_logic;			
			hps_io_hps_io_sdio_inst_CMD			: inout std_logic;
			hps_io_hps_io_sdio_inst_D0				: inout std_logic;
			hps_io_hps_io_sdio_inst_D1				: inout std_logic;
			hps_io_hps_io_sdio_inst_D2				: inout std_logic;
			hps_io_hps_io_sdio_inst_D3				: inout std_logic;

			hps_io_hps_io_usb1_inst_CLK			: in std_logic;
			hps_io_hps_io_usb1_inst_STP			: out std_logic;
			hps_io_hps_io_usb1_inst_DIR			: in std_logic;
			hps_io_hps_io_usb1_inst_NXT			: in std_logic;
			hps_io_hps_io_usb1_inst_D0				: inout std_logic;
			hps_io_hps_io_usb1_inst_D1				: inout std_logic;
			hps_io_hps_io_usb1_inst_D2				: inout std_logic;
			hps_io_hps_io_usb1_inst_D3				: inout std_logic;
			hps_io_hps_io_usb1_inst_D4				: inout std_logic;
			hps_io_hps_io_usb1_inst_D5				: inout std_logic;
			hps_io_hps_io_usb1_inst_D6				: inout std_logic;
			hps_io_hps_io_usb1_inst_D7				: inout std_logic;
			
			hps_io_hps_io_uart0_inst_RX			: in std_logic;
			hps_io_hps_io_uart0_inst_TX			: out std_logic;
			
			led_external_connection_export		: out std_logic_vector(9 downto 0);
			
			memory_mem_a								: out std_logic_vector(14 downto 0);
			memory_mem_ba								: out std_logic_vector(2 downto 0);			
			memory_mem_ck								: out std_logic;
			memory_mem_ck_n							: out std_logic;
			memory_mem_cke								: out std_logic;
			memory_mem_cs_n							: out std_logic;
			memory_mem_ras_n							: out std_logic;
			memory_mem_cas_n							: out std_logic;
			memory_mem_we_n							: out std_logic;
			memory_mem_reset_n						: out std_logic;
			memory_mem_dq								: inout std_logic_vector(31 downto 0);
			memory_mem_dqs								: inout std_logic_vector(3 downto 0);
			memory_mem_dqs_n							: inout std_logic_vector(3 downto 0);
			memory_mem_odt								: out std_logic;
			memory_mem_dm								: out std_logic_vector(3 downto 0);
			
			memory_oct_rzqin							: in std_logic;
			
			sdram_addr									: out std_logic_vector(10 downto 0);
			sdram_ba										: out std_logic_vector(1 downto 0);
			sdram_cas_n									: out std_logic;
			sdram_cke									: out std_logic;
			sdram_cs_n									: out std_logic;
			sdram_dq										: inout std_logic_vector(15 downto 0);
			sdram_dqm									: out std_logic_vector(1 downto 0);
			sdram_ras_n									: out std_logic;
			sdram_we_n									: out std_logic
		);
	end component arm_one_nios;
	
signal HPS_H2F_RST	: std_logic;
	
begin

	u0 : component arm_one_nios
		port map (
			clk_clk                         => CLOCK_50,
			reset_reset_n                   => '1',
			
			hps_0_h2f_reset_reset_n         => HPS_H2F_RST, 

			hps_io_hps_io_emac1_inst_TX_CLK => HPS_ENET_TX_CLK,
			hps_io_hps_io_emac1_inst_TX_CTL => HPS_ENET_TX_EN,
			hps_io_hps_io_emac1_inst_TXD0   => HPS_ENET_TX_DATA(0),
			hps_io_hps_io_emac1_inst_TXD1   => HPS_ENET_TX_DATA(1),
			hps_io_hps_io_emac1_inst_TXD2   => HPS_ENET_TX_DATA(2),
			hps_io_hps_io_emac1_inst_TXD3   => HPS_ENET_TX_DATA(3),
			hps_io_hps_io_emac1_inst_RX_CLK => HPS_ENET_RX_CLK,
			hps_io_hps_io_emac1_inst_RX_CTL => HPS_ENET_RX_DV,			
			hps_io_hps_io_emac1_inst_RXD0   => HPS_ENET_RX_DATA(0),
			hps_io_hps_io_emac1_inst_RXD1   => HPS_ENET_RX_DATA(1),
			hps_io_hps_io_emac1_inst_RXD2   => HPS_ENET_RX_DATA(2),
			hps_io_hps_io_emac1_inst_RXD3   => HPS_ENET_RX_DATA(3),
			hps_io_hps_io_emac1_inst_MDIO   => HPS_ENET_MDIO,
			hps_io_hps_io_emac1_inst_MDC    => HPS_ENET_MDC,
			
			hps_io_hps_io_sdio_inst_CLK     => HPS_SD_CLK,
			hps_io_hps_io_sdio_inst_CMD     => HPS_SD_CMD,
			hps_io_hps_io_sdio_inst_D0      => HPS_SD_DATA(0),
			hps_io_hps_io_sdio_inst_D1      => HPS_SD_DATA(1),
			hps_io_hps_io_sdio_inst_D2      => HPS_SD_DATA(2),
			hps_io_hps_io_sdio_inst_D3      => HPS_SD_DATA(3),
			
			hps_io_hps_io_usb1_inst_CLK     => HPS_USB_CLKOUT,
			hps_io_hps_io_usb1_inst_STP     => HPS_USB_STP,
			hps_io_hps_io_usb1_inst_DIR     => HPS_USB_DIR,
			hps_io_hps_io_usb1_inst_NXT     => HPS_USB_NXT,
			hps_io_hps_io_usb1_inst_D0      => HPS_USB_DATA(0),
			hps_io_hps_io_usb1_inst_D1      => HPS_USB_DATA(1),
			hps_io_hps_io_usb1_inst_D2      => HPS_USB_DATA(2),
			hps_io_hps_io_usb1_inst_D3      => HPS_USB_DATA(3),
			hps_io_hps_io_usb1_inst_D4      => HPS_USB_DATA(4),
			hps_io_hps_io_usb1_inst_D5      => HPS_USB_DATA(5),
			hps_io_hps_io_usb1_inst_D6      => HPS_USB_DATA(6),
			hps_io_hps_io_usb1_inst_D7      => HPS_USB_DATA(7),

			hps_io_hps_io_uart0_inst_RX     => HPS_UART_RX,
			hps_io_hps_io_uart0_inst_TX     => HPS_UART_TX,
			
			led_external_connection_export  => LEDR,
			
			memory_mem_a                    => HPS_DDR3_ADDR,
			memory_mem_ba                   => HPS_DDR3_BA,
			memory_mem_ck                   => HPS_DDR3_CK_P,
			memory_mem_ck_n                 => HPS_DDR3_CK_N,
			memory_mem_cke                  => HPS_DDR3_CKE,
			memory_mem_cs_n                 => HPS_DDR3_CS_N,
			memory_mem_ras_n                => HPS_DDR3_RAS_N,
			memory_mem_cas_n                => HPS_DDR3_CAS_N,
			memory_mem_we_n                 => HPS_DDR3_WE_N,
			memory_mem_reset_n              => HPS_DDR3_RESET_N,
			memory_mem_dq                   => HPS_DDR3_DQ,
			memory_mem_dqs                  => HPS_DDR3_DQS_P,
			memory_mem_dqs_n                => HPS_DDR3_DQS_N,
			memory_mem_odt                  => HPS_DDR3_ODT,
			memory_mem_dm                   => HPS_DDR3_DM,
			memory_oct_rzqin                => HPS_DDR3_RZQ,

			sdram_addr                      => SDRAM_ADDR,
			sdram_ba                        => SDRAM_BA,
			sdram_cas_n                     => SDRAM_CAS_N,
			sdram_cke                       => SDRAM_CKE,
			sdram_cs_n                      => SDRAM_CS_N,
			sdram_dq                        => SDRAM_DQ,
			sdram_dqm                       => SDRAM_DQM,
			sdram_ras_n                     => SDRAM_RAS_N,
			sdram_we_n                      => SDRAM_WE_N
		);
		
end main;
			
			
		
		
		
		
		
		
